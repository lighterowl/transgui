TranslationLanguage=Svenska

"Remote to local path mappings.~Examples:~/share=\\pch\share~/var/downloads/music=Z:\music"="Mappning fjärr- till lokala sökvägar.~Till exempel:~/share=\\pch\share~/var/downloads/musik=Z:\musik"
%d torrents=%d torrents
%d x %s (have %d)=%d x %s (har %d)
%dd=%dd
%dh=%dh
%dm=%dm
%ds=%ds
%s (%d hashfails)=%s (%d hashfel)
%s (%s done)=%s (%s klar)
%s downloaded=%s nedladdat
%s of %s downloaded=%s av %s nedladdat
%s%s%d downloading, %d seeding%s%s, %s=%s%s%d laddar ner, %d delar%s%s, %s
&Add torrent=Lägg till torrent
&All=&Alla
&Close=&Stäng
&Help=&Hjälp
&Ignore=&Ignorera
&No=&Nej
&OK=&OK
&Open=&Öppna
&Retry=&Försök igen
&Save=&Spara
&Torrent=Torrent
&Unlock=Lås upp
&Verify=Verifiera
&Yes=&Ja
'%s' has finished downloading='%s' är klar med nedladdningen
/s=/s
A new version of %s is available.~Your current version: %s~The new version: %s~Do you wish to open the Downloads web page?=A new version of %s is available.~Your current version: %s~The new version: %s~Do you wish to open the Downloads web page?
Abort=Avbryt
About=Om
Access violation=Åtkomstfel
Active time=Aktiv tid
Active=Aktiv
Add .part extension to incomplete files=Lägg till .part på ofullständiga filer
Add new torrent=Lägg till ny torrent
Add torrent link=Lägg till en torrentlänk
Add torrent=Lägg till torrent
Add tracker=Lägg till tracker
Added on=Lades till
Advanced=Avancerad
All torrents=Alla torrents
Allow encryption=Tillåt kryptering
Alternate bandwidth settings=Alternativa bandbreddsinställingar
Always auto-reconnect=Återanslut alltid automatiskt
Application Options (Ctrl+F9)=Applikationsinställningar (Ctrl+F9)
Application options=Programalternativ
Apply alternate bandwidth settings automatically=Använd alternativa bandbreddsinställningar automatiskt
Are you sure to delete connection '%s'?=Är du säker på att du vill ta bort anslutningen '%s'?
Are you sure to remove %d selected torrents and all their associated DATA?=är du säker på att du önskar att ta bort %d valda torrenter och alla tilhörande data?
Are you sure to remove %d selected torrents?=är du säker på att du önskar att ta bort %d valda torrenter?
Are you sure to remove torrent '%s' and all associated DATA?=Är du säker på att du vill ta bort '%s' och all tillhörande data?
Are you sure to remove torrent '%s'?=Är du säker på att du vill ta bort torrenten '%s'?
Are you sure to remove tracker '%s'?=Är du säker på att du vill ta bort trackern '%s'?
Ask for password=Fråga efter lösenord
Authentication required=Autentisering krävs
Authentication=Autentisering
Automatically add torrent links from the clipboard=Lägg automatiskt till torrent-länkar från urklipp
Average out transfer speeds to eliminate fluctuations=Jämna ut överföringshastigheten för att ta bort fluktuationer
average=genomsnitt
b=b
Bandwidth=Bandbredd
Browse=Bläddra
Cancel=Avbryt
Check for new version every=Sök efter nya versioner varje
Check for updates=Sök efter uppdateringar
Client=Klient
Close to tray=Stäng till aktivitetsfältet
Columns setup=Kolumninställning
Comment=Kommentar
Completed on=Avslutad den
Completed=Avslutad
Confirmation=Bekräftelse
Connect to %s=Anslut till %s
Connect to Transmission using proxy server=Anslut till Transmission via en proxyserver
Connect to Transmission=Anslut till Transmission
connected=ansluten
Connecting to daemon=Ansluter till server
Connection error occurred=Anslutningsfel har inträffat
Connection name=Namn på anslutningen
Connection refused=Anslutning avvisad
Connection timed out=Anslutningstidsavbrott
Consider active torrents as stalled when idle for=Anse att aktiva torrents är inaktiva efter
Copy file path to clipboard=Kopiera sökvägen till urklipp
Copy Magnet Link(s)=Kopiera magnetlänk(ar)
Copy=Kopiera
Could not connect to tracker==Kunde inte ansluta till tracker
Country=Land
Created on=Skapad
Cumulative=Kumulativ
Current=Aktuell
D: %s/s=D: %s/s
Data display=Datavisning
Data refresh interval when minimized=Uppdateringsintervall av data vid minimerad
Data refresh interval=Uppdateringsintervall av data
Days=Dagar
days=dagar
Default download folder on remote host=Nedladdningskatalog på Transmission-servern
Default=Standard
Delete a .torrent file after a successful addition=Ta bort .torrent-filen efter den lagts till
Delete destination folder=Ta bort destinationsmapp
Delete=Ta bort
Destination folder=Destinationsmapp
Development site=Webbplats för utveckling
Directory for incomplete files=Mapp för ofullständiga filer
Disconnect from Transmission=Stäng anslutningen till Transmission
Disconnected=Frånkopplad
Disk cache size=Storlek på diskcachen
Do you wish to enable automatic checking for a new version of %s?=Vill du aktivera automatisk kontroll av nya versioner av %s?
Don't download=Ladda inte ner
Donate to support further development=Donera för att stödja fortsatt utveckling
Donate via PayPal,WebMoney,Credit card=Donera via PayPal,WebMoney,Credit card
Donate!=Donera!
Done: %s=Klart: %s
Done=Färdig
Down limit=Nedladdningsgräns
Down speed=Nedladdningshastighet
Down=Ner
Download complete=Nedladdning klar
Download queue size=Storlek på nedladdningskön
Download speed=Nedladdingshastighet
Download speeds (KB/s)=Nedladdingshastighet (KB/s)
Download=Ladda ner
Downloaded=Nedladdad
Downloading torrent file=Laddar ner torrentfil
Downloading=Laddar ner
E&xit=Avsluta
Edit tracker=Redigera tracker
Enable blocklist=Aktivera blockeringslistan
Enable DHT=Aktivera DHT
Enable Local Peer Discovery=Aktivera Lokal Peer-upptäckt
Enable Peer Exchange=Aktivera Peer Exchange
Enable port forwarding=Aktivera portvidarebefordran
Enable µTP=Aktivera µTP
Encryption=Kryptering
Error checking for new version=Fel vid koll efter ny version
Error=Fel
ETA=ETA
Export settings=Exportera inställningar
File name=Filnamn
Files added=Filer tillagda
Files=Filer
Filter pane=Filterpanel
Finished=Färdig
Flag images archive is needed to display country flags.~Download this archive now?=Ett arkiv med flaggbilder är nödvändigt för att visa landsflaggor.~Vill du ladda ner denna nu?
Flags=Flaggor
Folder grouping=Gruppering av mappar
Font size=Storlek på typsnittet
for example: *.avi *.mkv=till exempel: *.avi *.mkv
Force start=Tvångsstarta
Free disk space=Ledigt diskutrymme
Free: %s=Ledigt: %s
From=Från
GB=GB
General=Allmänt
Geo IP database is needed to resolve country by IP address.~Download this database now?=En geo-IP databas är nödvändig för att visa vilket land en IP-adress tillhör.~Önskar du att ladda ner denna databasen nu??
Global bandwidth settings=Global bredbands inställningar
Global peer limit=Max antal globala kamrater
Global statistics=Global statistik
Handle .torrent files by %s=Hantera .torrent-filer via %s
Handle magnet links by %s=Hantera magnetlänkar via %s
Hash=Hash
Have=Har
Hide=Dölj
High priority=Hög prioritet
high=hög
Home page=Hemsida
Host not found=Värden kunde inte hittas
Host=Värd
ID=ID
Import settings=Importera inställningar
in swarm=i svärm
Inactive=Inaktiv
Incoming port is closed. Check your firewall settings=Inkommande port är stängd. Kontrollera brandväggs inställningarna
Incoming port tested successfully=Inkommande port är öppen
Incoming port=Inkommande port
Info pane=Informationspanel
Information=Information
Invalid name specified=Felaktigt namn angivet
KB/s=KB/s
KB=KB
Language=Språk
Last active=Senast aktiv
Left->Right=Vänster->Höger
License=Licens
Low priority=Låg prioritet
low=låg
Magnet Link=Magnetlänk
Manage connections to Transmission=Hantera anslutningar till Transmission
Manage connections=Hantera anslutningar
Max peers=Max antal peers
Maximum download speed=Max nedladdningshastighet
Maximum upload speed=Max uppladdningshastighet
MB=MB
Menu=Meny
Minimize to tray=Minimera till aktivitetsfältet
minutes=minuter
Misc=Diverse
Modify trackers=Ändra trackers
Move bottom=Flytta till botten av kön
Move down queue=Flytta ner i kön
Move down=Flytta ner
Move top=Flytta längst upp
Move torrent data from current location to new location=Flytta data från nuvarande plats till en ny plats
Move up queue=Flytta till toppen av kön
Move up=Flytta upp
Name=Namn
Network (WAN)=Nätverk (WAN)
New connection to Transmission=Ny anslutning till Transmission
New connection=Ny anslutning
New location for torrent data=Ny plats för torrent data
New=Ny
No host name specified=Inget värdnamn specifierat
No link was specified=Ingen länk specifierad
No proxy server specified=Ingen proxyserver specifierad
No to all=Nej till alla
No torrent location was specified=Ingen torrentplats var specifierad
No tracker URL was specified=Ingen trackeradress var specifierad
No tracker=Ingen tracker
No updates have been found.~You are running the latest version of %s=Inga uppdateringar hittades.~Du kör senaste versionen av %s
Normal priority=Normal prioritet
normal=normal
of=av
Open containing folder=Öppna målmapp
Open=Öppna
Other Winsock error=Annat Winsock-fel
Password=Lösenord
Path=Sökväg
Paths=Sökvägar
Peer limit=Peer begränsning
Peers=Peers
Pick random port on Transmission launch=Använd slumpad port när Transmission startar
Pieces=Delar
Please enter a password to connect to %s=Ange ett lösenord för att ansluta till %s
Please specify how %s will connect to a remote host running Transmission daemon (service)=Ange hur %s kommer ansluta till maskinen som kör Transmission-servern (service)
Port=Port
Prefer encryption=Föredra kryptering
Priority=Prioritet
Prompt for download options when adding a new torrent=Fråga om nedladdningsalternativ när en ny torrent läggs till
Properties=Egenskaper
Proxy password=Proxylösenord
Proxy port=Proxyport
Proxy server=Proxyserver
Proxy user name=Proxyanvändarnamn
Proxy=Proxy
Queue position=Köposition
Queue=Kö
Ratio=Förhållande
Reannounce (get more peers)=Tillkännage (skaffa flera peers)
Reconnect in %d seconds=Anslut på nytt om %d sekunder
Remaining: %s=Kvarvarande: %s
Remaining=Återstående
Remote host=Fjärrserver
Remove torrent and Data=Ta bort torrent och data
Remove torrent=Ta bort torrent
Remove tracker=Ta bort tracker
Remove=Ta bort
Rename=Byt namn
Require encryption=Kräv kryptering
Resolve country=Check land
Resolve host name=Check värdnamn
Right->Left (No Align)=Höger->Vänster (ingen centrering)
Right->Left (Reading Only)=Höger->Vänster (endast läsning)
Right->Left=Höger->Vänster
RPC path=RPC-sökväg
Save as=Spara som
seconds=sekunder
Seed ratio=Delningsförhållande
Seeding time=Uppladdningstid
Seeding=Delar
Seeds=Delare
Select a .torrent to open=Välj en .torrent att öppna
Select a folder for download=Välj nedladdningsmapp
Select all=Välj alla
Select none=Välj ingen
Select torrent location=Välj torrentplats
Selected: %s=Valt: %s
Set data location=Sätt dataplats
Setup columns=Ställ in kolumner
Share ratio=Delningsförhållande
Show advanced options=Visa avancerade alternativ
Show country flag=Visa flagga
Show notifications in tray icon=Visa notifieringar i ikonen i aktivitetsfältet
Show=Visa
Size left=Storlek kvar
Size to download=Storlek på nedladdning
Size=Storlek
skip=hoppa över
Speed limit menu items=Hastighetsbegränsningar
Start all torrents=Starta alla torrents
Start torrent=Starta torrent
Start=Starta
Statistics=Statistik
Status bar - Sizes=Statusrad - Storlekar
Status bar=Statusrad
Status=Status
Stop all torrents=Stoppa alla torrents
Stop all=Stoppa alla
Stop seeding when inactive for=Avsluta delning när inaktiv i
Stop torrent=Stoppa torrent
Stop=Stoppa
Stopped=Stoppad
System integration=Systemintegration
T&ools=Verktyg
TB=TB
Template:=Mall:
Test port=Testa porten
The block list has been updated successfully.~The list entries count: %d=Blockeringslistan blev uppdaterad.~Det är %d registrerade i listan
The directory for incomplete files was not specified=Mappen för ofullständiga filer var inte specifierad
The downloads directory was not specified=Nedladdningsmappen var inte specificerad
The invalid time value was entered=Ett ogiltig tidsvärde angavs
The maximum history of directories for storage of torrents=Maximal historik över mappar för torrentlagring
to=till
Toolbar=Verktygsfält
Torrent already exists in the list=Torrenten finns redan i listan
Torrent contents=Innehåll i torrent
Torrent data location=Dataplats for torrent
Torrent not registered with this tracker==Torrenten är inte registrerad hos denna tracker
Torrent properties=Egenskaper för torrent
Torrent verification may take a long time.~Are you sure to start verification of torrent '%s'?=Torrentverifikation kan ta lång tid.~Är du säker på att du vill starta torrentverifikation '%s'?
Torrent=Torrent
Torrents (*.torrent)|*.torrent|All files (*.*)|*.*=Torrenter (*.torrent)|*.torrent|Alla filar (*.*)|*.*
Torrents that are idle for N minuets aren't counted toward the Download queue or Upload queue=Torrents som är inaktiva under N minuter räknas inte mot Download kön eller Upload kön
Torrents verification may take a long time.~Are you sure to start verification of %d torrents?=Dataverifiering kan ta lång tid.~Är du säker på att du önskar att verifiera %d torrenter?
Torrents=Torrents
Total size=Total storlek
Total: %s=Totalt: %s
Tracker announce URL=Trackerns annonseringsadress
Tracker grouping=Trackergruppering
Tracker properties=Trackerinställningar
Tracker status=Trackerstatus
Tracker update on=Tracker uppdaterad den
Tracker=Tracker
Trackers=Trackers
Transfer=Överföring
Transmission options=Alternativ för Transmission
Transmission%s at %s:%s=Transmission%s på %s:%s
Tray icon always visible=Ikon i aktivitetsfältet alltid synlig
Tray icon=Ikon i aktivitetsfältet
U: %s/s=U: %s/s
Unable to execute "%s"=Kunde inte köra "%s"
Unable to extract flag image=Kunde inte hämta flaggbild
Unable to find path mapping.~Use the application's options to setup path mappings=Hittar inte katalogen.~Använd inställningarna under alternativ för detta programmet för att justera katalogen (path)
Unable to get files list=Kunde inte hämta fillista
Unable to load OpenSSL library files: %s and %s=Klarade inte att ladda OpenSSL biblioteks filerna: %s och %s från OpenSSL
Unauthorized User=Obehörig användare
Unknown=Okänt
Unlimited=Obegränsat
Up limit=Uppladdningsgräns
Up speed=Uppladdningshastighet
Up=Upp
Update blocklist=Uppdatera blockeringslista
Update complete=Uppdatering genomförd
Update GeoIP database=Uppdatera GeoIP-databas
Update in=Uppdaterar om
Update trackers for the existing torrent?=Uppdatera trackers för den existerande torrenten?
Updating=Uppdaterar
Upload queue size=Storlek på uppladdningskön
Upload speed=Uppladdningshastighet
Upload speeds (KB/s)=Uppladdningshastighet (KB/s)
Uploaded=Uppladdat
URL of a .torrent file or a magnet link=Adressen till en .torrent-fil eller en magnet-länk
Use alternate bandwidth settings=Använd alternativa bandbreddsinställningar
Use SSL=Använd SSL
User Menu=Användarmeny
User name=Användarnamn
Verify torrent=Verifiera torrents
Verifying=Verifierar
Version %s=Version %s
View=Visa
Visit home page=Besök hemsidan
Waiting=Väntar
Warning=Varning
Wasted=Bortkastat
Working=Arbetar
Yes to &All=Ja till &allt
You need to restart the application to apply changes=Du måste starta om programmet för att verkställa ändringarna
